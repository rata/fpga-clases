`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:44:48 10/01/2014 
// Design Name: 
// Module Name:    asd 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////



module asd(
output wire a,
input wire DO,
input wire DI,
input wire [5:0] RDADDR,
input wire RDCLK,
input wire REGCE,
input wire RST,
input wire WE,
input wire RDEN,
input wire [5:0] WRADDR,
input wire WRCLK,
input wire WREN
);

   BRAM_SDP_MACRO #(
      .BRAM_SIZE("18Kb"), // Target BRAM, "9Kb" or "18Kb" 
      .DEVICE("SPARTAN6"), // Target device: "VIRTEX5", "VIRTEX6", "SPARTAN6" 
      .WRITE_WIDTH(1),    // Valid values are 1-36
      .READ_WIDTH(1),     // Valid values are 1-36
      .DO_REG(0),         // Optional output register (0 or 1)
      .INIT_FILE ("NONE"),
      .SIM_COLLISION_CHECK ("ALL"), // Collision check enable "ALL", "WARNING_ONLY", 
                                    //   "GENERATE_X_ONLY" or "NONE" 
      .SRVAL(72'h000000000000000000), // Set/Reset value for port output
      .INIT(72'h000000000000000000),  // Initial values on output port
 //     .INIT_00(256'h00000000000000000000000000000000000000000000000000000000ffffffff),
      .INIT_00(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_01(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_02(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_03(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_04(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_05(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_06(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_07(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_08(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_09(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_0A(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_0B(256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
            
      // The next set of INIT_xx are for "18Kb" configuration only
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_30(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_31(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_32(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_33(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_34(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_35(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_36(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_37(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_38(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_39(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_3F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      
      // The next set of INITP_xx are for the parity bits
      .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
            
      // The next set of INITP_xx are for "18Kb" configuration only
      .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000)
   )

BRAM_SDP_MACRO_inst (
      .DO(DO),         // Output read data port, width defined by READ_WIDTH parameter
      .DI(DI),         // Input write data port, width defined by WRITE_WIDTH parameter
      .RDADDR(RDADDR), // Input read address, width defined by read port depth
      .RDCLK(RDCLK),   // 1-bit input read clock
      .RDEN(RDEN),     // 1-bit input read port enable
      .REGCE(REGCE),   // 1-bit input read output register enable
      .RST(RST),       // 1-bit input reset      
      .WE(WE),         // Input write enable, width defined by write port depth
      .WRADDR(WRADDR), // Input write address, width defined by write port depth
      .WRCLK(WRCLK),   // 1-bit input write clock
      .WREN(WREN)      // 1-bit input write port enable
   );

assign a = DO;
endmodule 
